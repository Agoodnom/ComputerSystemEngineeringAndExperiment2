`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/10/09 23:52:41
// Design Name: 
// Module Name: 1_bit_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module one_bit_tb;

reg in_a,in_b;
wire out_c,out_d,out_e,out_f;

one_bit sim(
.a(in_a),
.b(in_b),
.c(out_c),
.d(out_d),
.e(out_e),
.f(out_f)
);

initial
begin
    in_a = 1'b0;
    in_b = 1'b0;
end

always@(in_a or in_b)
begin
    in_a <=#4 ~in_a;
    in_b <=#2 ~in_b;
end
endmodule
